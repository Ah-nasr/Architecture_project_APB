library verilog;
use verilog.vl_types.all;
entity master_bridge_tb is
end master_bridge_tb;
